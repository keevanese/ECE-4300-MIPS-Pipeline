`timescale 1ns / 1ps
/*
ALU: performs arithmetic and logic operations based on 3-bit control.
*/

module alu(
    input  wire [31:0] a,       // source register
    input  wire [31:0] b,       // second operand
    input  wire [2:0]  control, // from alu_control
    output reg  [31:0] result,
    output wire        zero
);

    // Must match alu_control encodings
    localparam ALU_ADD = 3'b010;
    localparam ALU_SUB = 3'b110;
    localparam ALU_AND = 3'b000;
    localparam ALU_OR  = 3'b001;
    localparam ALU_SLT = 3'b111;

    initial result = 32'd0;

    always @* begin
        case (control)
            ALU_ADD: result = a + b;
            ALU_SUB: result = a - b;
            ALU_AND: result = a & b;
            ALU_OR : result = a | b;
            ALU_SLT: result = ($signed(a) < $signed(b)) ? 32'd1 : 32'd0;
            default: result = 32'hXXXXXXXX;
        endcase
    end

    // zero flag: 1 if result == 0
    assign zero = (result == 32'd0);

endmodule